module VexRiscv(
 input      [31:0]   externalResetVector,
  input               timerInterrupt,
  input               softwareInterrupt,
  input      [31:0]   externalInterruptArray,
  output              debug_resetOut,
  output              iBusAxi_ar_valid,
  input               iBusAxi_ar_ready,
  output     [31:0]   iBusAxi_ar_payload_addr,
  output     [0:0]    iBusAxi_ar_payload_id,
  output     [3:0]    iBusAxi_ar_payload_region,
  output     [7:0]    iBusAxi_ar_payload_len,
  output     [2:0]    iBusAxi_ar_payload_size,
  output     [1:0]    iBusAxi_ar_payload_burst,
  output     [0:0]    iBusAxi_ar_payload_lock,
  output     [3:0]    iBusAxi_ar_payload_cache,
  output     [3:0]    iBusAxi_ar_payload_qos,
  output     [2:0]    iBusAxi_ar_payload_prot,
  input               iBusAxi_r_valid,
  output              iBusAxi_r_ready,
  input      [31:0]   iBusAxi_r_payload_data,
  input      [0:0]    iBusAxi_r_payload_id,
  input      [1:0]    iBusAxi_r_payload_resp,
  input               iBusAxi_r_payload_last,
  output              dBusAxi_aw_valid,
  input               dBusAxi_aw_ready,
  output     [31:0]   dBusAxi_aw_payload_addr,
  output     [0:0]    dBusAxi_aw_payload_id,
  output     [3:0]    dBusAxi_aw_payload_region,
  output     [7:0]    dBusAxi_aw_payload_len,
  output     [2:0]    dBusAxi_aw_payload_size,
  output     [1:0]    dBusAxi_aw_payload_burst,
  output     [0:0]    dBusAxi_aw_payload_lock,
  output     [3:0]    dBusAxi_aw_payload_cache,
  output     [3:0]    dBusAxi_aw_payload_qos,
  output     [2:0]    dBusAxi_aw_payload_prot,
  output              dBusAxi_w_valid,
  input               dBusAxi_w_ready,
  output     [31:0]   dBusAxi_w_payload_data,
  output     [3:0]    dBusAxi_w_payload_strb,
  output              dBusAxi_w_payload_last,
  input               dBusAxi_b_valid,
  output              dBusAxi_b_ready,
  input      [0:0]    dBusAxi_b_payload_id,
  input      [1:0]    dBusAxi_b_payload_resp,
  output              dBusAxi_ar_valid,
  input               dBusAxi_ar_ready,
  output     [31:0]   dBusAxi_ar_payload_addr,
  output     [0:0]    dBusAxi_ar_payload_id,
  output     [3:0]    dBusAxi_ar_payload_region,
  output     [7:0]    dBusAxi_ar_payload_len,
  output     [2:0]    dBusAxi_ar_payload_size,
  output     [1:0]    dBusAxi_ar_payload_burst,
  output     [0:0]    dBusAxi_ar_payload_lock,
  output     [3:0]    dBusAxi_ar_payload_cache,
  output     [3:0]    dBusAxi_ar_payload_qos,
  output     [2:0]    dBusAxi_ar_payload_prot,
  input               dBusAxi_r_valid,
  output              dBusAxi_r_ready,
  input      [31:0]   dBusAxi_r_payload_data,
  input      [0:0]    dBusAxi_r_payload_id,
  input      [1:0]    dBusAxi_r_payload_resp,
  input               dBusAxi_r_payload_last,
  input               jtag_tms,
  input               jtag_tdi,
  output              jtag_tdo,
  input               jtag_tck,
  input               clk,
  input               reset,
  input               debugReset
);

wire soc_basesoc_vexriscv_cfu_bus_cmd_valid;
wire soc_basesoc_vexriscv_cfu_bus_cmd_ready;
wire [9:0] soc_basesoc_vexriscv_cfu_bus_cmd_payload_function_id;
wire [31:0] soc_basesoc_vexriscv_cfu_bus_cmd_payload_inputs_0;
wire [31:0] soc_basesoc_vexriscv_cfu_bus_cmd_payload_inputs_1;
wire soc_basesoc_vexriscv_cfu_bus_rsp_valid;
wire soc_basesoc_vexriscv_cfu_bus_rsp_ready;
wire [31:0] soc_basesoc_vexriscv_cfu_bus_rsp_payload_outputs_0;
//reg  [31:0] soc_basesoc_vexriscv = 32'd0;

Cfu Cfu(
	.clk(clk),
	.cmd_payload_function_id(soc_basesoc_vexriscv_cfu_bus_cmd_payload_function_id),
	.cmd_payload_inputs_0(soc_basesoc_vexriscv_cfu_bus_cmd_payload_inputs_0),
	.cmd_payload_inputs_1(soc_basesoc_vexriscv_cfu_bus_cmd_payload_inputs_1),
	.cmd_valid(soc_basesoc_vexriscv_cfu_bus_cmd_valid),
	.reset(reset),
	.rsp_ready(soc_basesoc_vexriscv_cfu_bus_rsp_ready),
	.cmd_ready(soc_basesoc_vexriscv_cfu_bus_cmd_ready),
	.rsp_payload_outputs_0(soc_basesoc_vexriscv_cfu_bus_rsp_payload_outputs_0),
	.rsp_valid(soc_basesoc_vexriscv_cfu_bus_rsp_valid)
);


VexRiscv_FullCfu VexRiscv1(
	.CfuPlugin_bus_cmd_ready(soc_basesoc_vexriscv_cfu_bus_cmd_ready),
	.CfuPlugin_bus_rsp_payload_outputs_0(soc_basesoc_vexriscv_cfu_bus_rsp_payload_outputs_0),
	.CfuPlugin_bus_rsp_valid(soc_basesoc_vexriscv_cfu_bus_rsp_valid),
	.CfuPlugin_bus_cmd_payload_function_id(soc_basesoc_vexriscv_cfu_bus_cmd_payload_function_id),
	.CfuPlugin_bus_cmd_payload_inputs_0(soc_basesoc_vexriscv_cfu_bus_cmd_payload_inputs_0),
	.CfuPlugin_bus_cmd_payload_inputs_1(soc_basesoc_vexriscv_cfu_bus_cmd_payload_inputs_1),
	.CfuPlugin_bus_cmd_valid(soc_basesoc_vexriscv_cfu_bus_cmd_valid),
	.CfuPlugin_bus_rsp_ready(soc_basesoc_vexriscv_cfu_bus_rsp_ready),
	.clk(clk),                            
	.reset(reset),      
    .dBusAxi_aw_valid(dBusAxi_aw_valid),      
    .dBusAxi_aw_ready(dBusAxi_aw_ready),      
    .dBusAxi_aw_payload_addr(dBusAxi_aw_payload_addr),       
    .dBusAxi_aw_payload_id(dBusAxi_aw_payload_id ),         
    .dBusAxi_aw_payload_region(dBusAxi_aw_payload_region),      
    .dBusAxi_aw_payload_len(dBusAxi_aw_payload_len),        
    .dBusAxi_aw_payload_size(dBusAxi_aw_payload_size),        
    .dBusAxi_aw_payload_burst(dBusAxi_aw_payload_burst),       
    .dBusAxi_aw_payload_lock(dBusAxi_aw_payload_lock),       
    .dBusAxi_aw_payload_cache(dBusAxi_aw_payload_cache),      
    .dBusAxi_aw_payload_qos(dBusAxi_aw_payload_qos),         
    .dBusAxi_aw_payload_prot(dBusAxi_aw_payload_prot),       
    .dBusAxi_w_valid(dBusAxi_w_valid),        
    .dBusAxi_w_ready(dBusAxi_w_ready),       
    .dBusAxi_w_payload_data(dBusAxi_w_payload_data),         
    .dBusAxi_w_payload_strb(dBusAxi_w_payload_strb),         
    .dBusAxi_w_payload_last(dBusAxi_w_payload_last),         
    .dBusAxi_b_valid(dBusAxi_b_valid),      
    .dBusAxi_b_ready(dBusAxi_b_ready),        
    .dBusAxi_b_payload_id(dBusAxi_b_payload_id),           
    .dBusAxi_b_payload_resp(dBusAxi_b_payload_resp),         
    .dBusAxi_ar_valid(dBusAxi_ar_valid),       
    .dBusAxi_ar_ready(dBusAxi_ar_ready),       
    .dBusAxi_ar_payload_addr(dBusAxi_ar_payload_addr),        
    .dBusAxi_ar_payload_id(dBusAxi_ar_payload_id),         
    .dBusAxi_ar_payload_region(dBusAxi_ar_payload_region),     
    .dBusAxi_ar_payload_len(dBusAxi_ar_payload_len),         
    .dBusAxi_ar_payload_size(dBusAxi_ar_payload_size),       
    .dBusAxi_ar_payload_burst(dBusAxi_ar_payload_burst),       
    .dBusAxi_ar_payload_lock(dBusAxi_ar_payload_lock),       
    .dBusAxi_ar_payload_cache(dBusAxi_ar_payload_cache),       
    .dBusAxi_ar_payload_qos(dBusAxi_ar_payload_qos),         
    .dBusAxi_ar_payload_prot(dBusAxi_ar_payload_prot),        
    .dBusAxi_r_valid(dBusAxi_r_valid),       
    .dBusAxi_r_ready(dBusAxi_r_ready),      
    .dBusAxi_r_payload_data(dBusAxi_r_payload_data),         
    .dBusAxi_r_payload_id(dBusAxi_r_payload_id),           
    .dBusAxi_r_payload_resp(dBusAxi_r_payload_resp),        
    .dBusAxi_r_payload_last(dBusAxi_r_payload_last),       
    .iBusAxi_ar_valid(iBusAxi_ar_valid),       
    .iBusAxi_ar_ready(iBusAxi_ar_ready),       
    .iBusAxi_ar_payload_addr(iBusAxi_ar_payload_addr),        
    .iBusAxi_ar_payload_id(iBusAxi_ar_payload_id),          
    .iBusAxi_ar_payload_region(iBusAxi_ar_payload_region),      
    .iBusAxi_ar_payload_len(iBusAxi_ar_payload_len),         
    .iBusAxi_ar_payload_size(iBusAxi_ar_payload_size),      
    .iBusAxi_ar_payload_burst(iBusAxi_ar_payload_burst),       
    .iBusAxi_ar_payload_lock(iBusAxi_ar_payload_lock),       
    .iBusAxi_ar_payload_cache(iBusAxi_ar_payload_cache),       
    .iBusAxi_ar_payload_qos(iBusAxi_ar_payload_qos),       
    .iBusAxi_ar_payload_prot(iBusAxi_ar_payload_prot),      
    .iBusAxi_r_valid(iBusAxi_r_valid),        
    .iBusAxi_r_ready(iBusAxi_r_ready),       
    .iBusAxi_r_payload_data(iBusAxi_r_payload_data),         
    .iBusAxi_r_payload_id(iBusAxi_r_payload_id),           
    .iBusAxi_r_payload_resp(iBusAxi_r_payload_resp),         
    .iBusAxi_r_payload_last(iBusAxi_r_payload_last),   
    .externalResetVector(externalResetVector),
    .timerInterrupt(timerInterrupt),
    .softwareInterrupt(softwareInterrupt),
     .externalInterruptArray(externalInterruptArray),
     .debug_resetOut(debug_resetOut),     
     .debugReset(debugReset),                 
	.jtag_tms(jtag_tms),                                    
	.jtag_tdi(jtag_tdi),                                     
	.jtag_tdo(jtag_tdo),                                    
	.jtag_tck(jtag_tck)                                      

);
endmodule
